// sopc4.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module sopc4 (
		input  wire       clk_clk,        //     clk.clk
		input  wire [7:0] in0_export,     //     in0.export
		input  wire [7:0] in1_export,     //     in1.export
		input  wire [7:0] in2_export,     //     in2.export
		input  wire [7:0] in3_export,     //     in3.export
		input  wire [7:0] in4_export,     //     in4.export
		input  wire [7:0] in5_export,     //     in5.export
		input  wire [7:0] in6_export,     //     in6.export
		input  wire [7:0] in7_export,     //     in7.export
		input  wire [7:0] in_aux_export,  //  in_aux.export
		output wire [7:0] out0_export,    //    out0.export
		output wire [7:0] out1_export,    //    out1.export
		output wire [7:0] out2_export,    //    out2.export
		output wire [7:0] out3_export,    //    out3.export
		output wire [7:0] out4_export,    //    out4.export
		output wire [7:0] out5_export,    //    out5.export
		output wire [7:0] out6_export,    //    out6.export
		output wire [7:0] out7_export,    //    out7.export
		output wire [7:0] out_aux_export, // out_aux.export
		input  wire       reset_reset_n   //   reset.reset_n
	);

	wire  [31:0] cpu_data_master_readdata;                             // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                          // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                          // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [19:0] cpu_data_master_address;                              // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                           // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                 // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                        // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                            // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                      // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                   // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [19:0] cpu_instruction_master_address;                       // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                          // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                 // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;    // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest; // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;       // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;        // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;       // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;    // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;    // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;        // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;           // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;     // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;          // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;      // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_memory_s1_chipselect;               // mm_interconnect_0:memory_s1_chipselect -> memory:chipselect
	wire  [31:0] mm_interconnect_0_memory_s1_readdata;                 // memory:readdata -> mm_interconnect_0:memory_s1_readdata
	wire  [15:0] mm_interconnect_0_memory_s1_address;                  // mm_interconnect_0:memory_s1_address -> memory:address
	wire   [3:0] mm_interconnect_0_memory_s1_byteenable;               // mm_interconnect_0:memory_s1_byteenable -> memory:byteenable
	wire         mm_interconnect_0_memory_s1_write;                    // mm_interconnect_0:memory_s1_write -> memory:write
	wire  [31:0] mm_interconnect_0_memory_s1_writedata;                // mm_interconnect_0:memory_s1_writedata -> memory:writedata
	wire         mm_interconnect_0_memory_s1_clken;                    // mm_interconnect_0:memory_s1_clken -> memory:clken
	wire  [31:0] mm_interconnect_0_in_aux_s1_readdata;                 // in_aux:readdata -> mm_interconnect_0:in_aux_s1_readdata
	wire   [1:0] mm_interconnect_0_in_aux_s1_address;                  // mm_interconnect_0:in_aux_s1_address -> in_aux:address
	wire         mm_interconnect_0_out_aux_s1_chipselect;              // mm_interconnect_0:out_aux_s1_chipselect -> out_aux:chipselect
	wire  [31:0] mm_interconnect_0_out_aux_s1_readdata;                // out_aux:readdata -> mm_interconnect_0:out_aux_s1_readdata
	wire   [1:0] mm_interconnect_0_out_aux_s1_address;                 // mm_interconnect_0:out_aux_s1_address -> out_aux:address
	wire         mm_interconnect_0_out_aux_s1_write;                   // mm_interconnect_0:out_aux_s1_write -> out_aux:write_n
	wire  [31:0] mm_interconnect_0_out_aux_s1_writedata;               // mm_interconnect_0:out_aux_s1_writedata -> out_aux:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                  // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                   // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                     // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                 // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire  [31:0] mm_interconnect_0_in7_s1_readdata;                    // in7:readdata -> mm_interconnect_0:in7_s1_readdata
	wire   [1:0] mm_interconnect_0_in7_s1_address;                     // mm_interconnect_0:in7_s1_address -> in7:address
	wire  [31:0] mm_interconnect_0_in6_s1_readdata;                    // in6:readdata -> mm_interconnect_0:in6_s1_readdata
	wire   [1:0] mm_interconnect_0_in6_s1_address;                     // mm_interconnect_0:in6_s1_address -> in6:address
	wire  [31:0] mm_interconnect_0_in5_s1_readdata;                    // in5:readdata -> mm_interconnect_0:in5_s1_readdata
	wire   [1:0] mm_interconnect_0_in5_s1_address;                     // mm_interconnect_0:in5_s1_address -> in5:address
	wire  [31:0] mm_interconnect_0_in4_s1_readdata;                    // in4:readdata -> mm_interconnect_0:in4_s1_readdata
	wire   [1:0] mm_interconnect_0_in4_s1_address;                     // mm_interconnect_0:in4_s1_address -> in4:address
	wire  [31:0] mm_interconnect_0_in3_s1_readdata;                    // in3:readdata -> mm_interconnect_0:in3_s1_readdata
	wire   [1:0] mm_interconnect_0_in3_s1_address;                     // mm_interconnect_0:in3_s1_address -> in3:address
	wire  [31:0] mm_interconnect_0_in2_s1_readdata;                    // in2:readdata -> mm_interconnect_0:in2_s1_readdata
	wire   [1:0] mm_interconnect_0_in2_s1_address;                     // mm_interconnect_0:in2_s1_address -> in2:address
	wire  [31:0] mm_interconnect_0_in1_s1_readdata;                    // in1:readdata -> mm_interconnect_0:in1_s1_readdata
	wire   [1:0] mm_interconnect_0_in1_s1_address;                     // mm_interconnect_0:in1_s1_address -> in1:address
	wire  [31:0] mm_interconnect_0_in0_s1_readdata;                    // in0:readdata -> mm_interconnect_0:in0_s1_readdata
	wire   [1:0] mm_interconnect_0_in0_s1_address;                     // mm_interconnect_0:in0_s1_address -> in0:address
	wire         mm_interconnect_0_out0_s1_chipselect;                 // mm_interconnect_0:out0_s1_chipselect -> out0:chipselect
	wire  [31:0] mm_interconnect_0_out0_s1_readdata;                   // out0:readdata -> mm_interconnect_0:out0_s1_readdata
	wire   [1:0] mm_interconnect_0_out0_s1_address;                    // mm_interconnect_0:out0_s1_address -> out0:address
	wire         mm_interconnect_0_out0_s1_write;                      // mm_interconnect_0:out0_s1_write -> out0:write_n
	wire  [31:0] mm_interconnect_0_out0_s1_writedata;                  // mm_interconnect_0:out0_s1_writedata -> out0:writedata
	wire         mm_interconnect_0_out1_s1_chipselect;                 // mm_interconnect_0:out1_s1_chipselect -> out1:chipselect
	wire  [31:0] mm_interconnect_0_out1_s1_readdata;                   // out1:readdata -> mm_interconnect_0:out1_s1_readdata
	wire   [1:0] mm_interconnect_0_out1_s1_address;                    // mm_interconnect_0:out1_s1_address -> out1:address
	wire         mm_interconnect_0_out1_s1_write;                      // mm_interconnect_0:out1_s1_write -> out1:write_n
	wire  [31:0] mm_interconnect_0_out1_s1_writedata;                  // mm_interconnect_0:out1_s1_writedata -> out1:writedata
	wire         mm_interconnect_0_out2_s1_chipselect;                 // mm_interconnect_0:out2_s1_chipselect -> out2:chipselect
	wire  [31:0] mm_interconnect_0_out2_s1_readdata;                   // out2:readdata -> mm_interconnect_0:out2_s1_readdata
	wire   [1:0] mm_interconnect_0_out2_s1_address;                    // mm_interconnect_0:out2_s1_address -> out2:address
	wire         mm_interconnect_0_out2_s1_write;                      // mm_interconnect_0:out2_s1_write -> out2:write_n
	wire  [31:0] mm_interconnect_0_out2_s1_writedata;                  // mm_interconnect_0:out2_s1_writedata -> out2:writedata
	wire         mm_interconnect_0_out3_s1_chipselect;                 // mm_interconnect_0:out3_s1_chipselect -> out3:chipselect
	wire  [31:0] mm_interconnect_0_out3_s1_readdata;                   // out3:readdata -> mm_interconnect_0:out3_s1_readdata
	wire   [1:0] mm_interconnect_0_out3_s1_address;                    // mm_interconnect_0:out3_s1_address -> out3:address
	wire         mm_interconnect_0_out3_s1_write;                      // mm_interconnect_0:out3_s1_write -> out3:write_n
	wire  [31:0] mm_interconnect_0_out3_s1_writedata;                  // mm_interconnect_0:out3_s1_writedata -> out3:writedata
	wire         mm_interconnect_0_out4_s1_chipselect;                 // mm_interconnect_0:out4_s1_chipselect -> out4:chipselect
	wire  [31:0] mm_interconnect_0_out4_s1_readdata;                   // out4:readdata -> mm_interconnect_0:out4_s1_readdata
	wire   [1:0] mm_interconnect_0_out4_s1_address;                    // mm_interconnect_0:out4_s1_address -> out4:address
	wire         mm_interconnect_0_out4_s1_write;                      // mm_interconnect_0:out4_s1_write -> out4:write_n
	wire  [31:0] mm_interconnect_0_out4_s1_writedata;                  // mm_interconnect_0:out4_s1_writedata -> out4:writedata
	wire         mm_interconnect_0_out5_s1_chipselect;                 // mm_interconnect_0:out5_s1_chipselect -> out5:chipselect
	wire  [31:0] mm_interconnect_0_out5_s1_readdata;                   // out5:readdata -> mm_interconnect_0:out5_s1_readdata
	wire   [1:0] mm_interconnect_0_out5_s1_address;                    // mm_interconnect_0:out5_s1_address -> out5:address
	wire         mm_interconnect_0_out5_s1_write;                      // mm_interconnect_0:out5_s1_write -> out5:write_n
	wire  [31:0] mm_interconnect_0_out5_s1_writedata;                  // mm_interconnect_0:out5_s1_writedata -> out5:writedata
	wire         mm_interconnect_0_out6_s1_chipselect;                 // mm_interconnect_0:out6_s1_chipselect -> out6:chipselect
	wire  [31:0] mm_interconnect_0_out6_s1_readdata;                   // out6:readdata -> mm_interconnect_0:out6_s1_readdata
	wire   [1:0] mm_interconnect_0_out6_s1_address;                    // mm_interconnect_0:out6_s1_address -> out6:address
	wire         mm_interconnect_0_out6_s1_write;                      // mm_interconnect_0:out6_s1_write -> out6:write_n
	wire  [31:0] mm_interconnect_0_out6_s1_writedata;                  // mm_interconnect_0:out6_s1_writedata -> out6:writedata
	wire         mm_interconnect_0_out7_s1_chipselect;                 // mm_interconnect_0:out7_s1_chipselect -> out7:chipselect
	wire  [31:0] mm_interconnect_0_out7_s1_readdata;                   // out7:readdata -> mm_interconnect_0:out7_s1_readdata
	wire   [1:0] mm_interconnect_0_out7_s1_address;                    // mm_interconnect_0:out7_s1_address -> out7:address
	wire         mm_interconnect_0_out7_s1_write;                      // mm_interconnect_0:out7_s1_write -> out7:write_n
	wire  [31:0] mm_interconnect_0_out7_s1_writedata;                  // mm_interconnect_0:out7_s1_writedata -> out7:writedata
	wire         irq_mapper_receiver0_irq;                             // jtag:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                             // timer:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_irq_irq;                                          // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [cpu:reset_n, in0:reset_n, in1:reset_n, in2:reset_n, in3:reset_n, in4:reset_n, in5:reset_n, in6:reset_n, in7:reset_n, in_aux:reset_n, irq_mapper:reset, jtag:rst_n, memory:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, out0:reset_n, out1:reset_n, out2:reset_n, out3:reset_n, out4:reset_n, out5:reset_n, out6:reset_n, out7:reset_n, out_aux:reset_n, rst_translator:in_reset, sysid:reset_n, timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                   // rst_controller:reset_req -> [cpu:reset_req, memory:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                        // cpu:debug_reset_request -> rst_controller:reset_in1

	sopc4_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	sopc4_in0 in0 (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_in0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in0_s1_readdata), //                    .readdata
		.in_port  (in0_export)                         // external_connection.export
	);

	sopc4_in0 in1 (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_in1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in1_s1_readdata), //                    .readdata
		.in_port  (in1_export)                         // external_connection.export
	);

	sopc4_in0 in2 (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_in2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in2_s1_readdata), //                    .readdata
		.in_port  (in2_export)                         // external_connection.export
	);

	sopc4_in0 in3 (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_in3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in3_s1_readdata), //                    .readdata
		.in_port  (in3_export)                         // external_connection.export
	);

	sopc4_in0 in4 (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_in4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in4_s1_readdata), //                    .readdata
		.in_port  (in4_export)                         // external_connection.export
	);

	sopc4_in0 in5 (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_in5_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in5_s1_readdata), //                    .readdata
		.in_port  (in5_export)                         // external_connection.export
	);

	sopc4_in0 in6 (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_in6_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in6_s1_readdata), //                    .readdata
		.in_port  (in6_export)                         // external_connection.export
	);

	sopc4_in0 in7 (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_in7_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in7_s1_readdata), //                    .readdata
		.in_port  (in7_export)                         // external_connection.export
	);

	sopc4_in0 in_aux (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_in_aux_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in_aux_s1_readdata), //                    .readdata
		.in_port  (in_aux_export)                         // external_connection.export
	);

	sopc4_jtag jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	sopc4_memory memory (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	sopc4_out0 out0 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_out0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out0_s1_readdata),   //                    .readdata
		.out_port   (out0_export)                           // external_connection.export
	);

	sopc4_out0 out1 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_out1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out1_s1_readdata),   //                    .readdata
		.out_port   (out1_export)                           // external_connection.export
	);

	sopc4_out0 out2 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_out2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out2_s1_readdata),   //                    .readdata
		.out_port   (out2_export)                           // external_connection.export
	);

	sopc4_out0 out3 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_out3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out3_s1_readdata),   //                    .readdata
		.out_port   (out3_export)                           // external_connection.export
	);

	sopc4_out0 out4 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_out4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out4_s1_readdata),   //                    .readdata
		.out_port   (out4_export)                           // external_connection.export
	);

	sopc4_out0 out5 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_out5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out5_s1_readdata),   //                    .readdata
		.out_port   (out5_export)                           // external_connection.export
	);

	sopc4_out0 out6 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_out6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out6_s1_readdata),   //                    .readdata
		.out_port   (out6_export)                           // external_connection.export
	);

	sopc4_out0 out7 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_out7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out7_s1_readdata),   //                    .readdata
		.out_port   (out7_export)                           // external_connection.export
	);

	sopc4_out0 out_aux (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_out_aux_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out_aux_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out_aux_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out_aux_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out_aux_s1_readdata),   //                    .readdata
		.out_port   (out_aux_export)                           // external_connection.export
	);

	sopc4_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	sopc4_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	sopc4_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                         (clk_clk),                                              //                       clk_0_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address               (cpu_data_master_address),                              //                 cpu_data_master.address
		.cpu_data_master_waitrequest           (cpu_data_master_waitrequest),                          //                                .waitrequest
		.cpu_data_master_byteenable            (cpu_data_master_byteenable),                           //                                .byteenable
		.cpu_data_master_read                  (cpu_data_master_read),                                 //                                .read
		.cpu_data_master_readdata              (cpu_data_master_readdata),                             //                                .readdata
		.cpu_data_master_readdatavalid         (cpu_data_master_readdatavalid),                        //                                .readdatavalid
		.cpu_data_master_write                 (cpu_data_master_write),                                //                                .write
		.cpu_data_master_writedata             (cpu_data_master_writedata),                            //                                .writedata
		.cpu_data_master_debugaccess           (cpu_data_master_debugaccess),                          //                                .debugaccess
		.cpu_instruction_master_address        (cpu_instruction_master_address),                       //          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest    (cpu_instruction_master_waitrequest),                   //                                .waitrequest
		.cpu_instruction_master_read           (cpu_instruction_master_read),                          //                                .read
		.cpu_instruction_master_readdata       (cpu_instruction_master_readdata),                      //                                .readdata
		.cpu_instruction_master_readdatavalid  (cpu_instruction_master_readdatavalid),                 //                                .readdatavalid
		.cpu_debug_mem_slave_address           (mm_interconnect_0_cpu_debug_mem_slave_address),        //             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write             (mm_interconnect_0_cpu_debug_mem_slave_write),          //                                .write
		.cpu_debug_mem_slave_read              (mm_interconnect_0_cpu_debug_mem_slave_read),           //                                .read
		.cpu_debug_mem_slave_readdata          (mm_interconnect_0_cpu_debug_mem_slave_readdata),       //                                .readdata
		.cpu_debug_mem_slave_writedata         (mm_interconnect_0_cpu_debug_mem_slave_writedata),      //                                .writedata
		.cpu_debug_mem_slave_byteenable        (mm_interconnect_0_cpu_debug_mem_slave_byteenable),     //                                .byteenable
		.cpu_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),    //                                .waitrequest
		.cpu_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),    //                                .debugaccess
		.in0_s1_address                        (mm_interconnect_0_in0_s1_address),                     //                          in0_s1.address
		.in0_s1_readdata                       (mm_interconnect_0_in0_s1_readdata),                    //                                .readdata
		.in1_s1_address                        (mm_interconnect_0_in1_s1_address),                     //                          in1_s1.address
		.in1_s1_readdata                       (mm_interconnect_0_in1_s1_readdata),                    //                                .readdata
		.in2_s1_address                        (mm_interconnect_0_in2_s1_address),                     //                          in2_s1.address
		.in2_s1_readdata                       (mm_interconnect_0_in2_s1_readdata),                    //                                .readdata
		.in3_s1_address                        (mm_interconnect_0_in3_s1_address),                     //                          in3_s1.address
		.in3_s1_readdata                       (mm_interconnect_0_in3_s1_readdata),                    //                                .readdata
		.in4_s1_address                        (mm_interconnect_0_in4_s1_address),                     //                          in4_s1.address
		.in4_s1_readdata                       (mm_interconnect_0_in4_s1_readdata),                    //                                .readdata
		.in5_s1_address                        (mm_interconnect_0_in5_s1_address),                     //                          in5_s1.address
		.in5_s1_readdata                       (mm_interconnect_0_in5_s1_readdata),                    //                                .readdata
		.in6_s1_address                        (mm_interconnect_0_in6_s1_address),                     //                          in6_s1.address
		.in6_s1_readdata                       (mm_interconnect_0_in6_s1_readdata),                    //                                .readdata
		.in7_s1_address                        (mm_interconnect_0_in7_s1_address),                     //                          in7_s1.address
		.in7_s1_readdata                       (mm_interconnect_0_in7_s1_readdata),                    //                                .readdata
		.in_aux_s1_address                     (mm_interconnect_0_in_aux_s1_address),                  //                       in_aux_s1.address
		.in_aux_s1_readdata                    (mm_interconnect_0_in_aux_s1_readdata),                 //                                .readdata
		.jtag_avalon_jtag_slave_address        (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //          jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write          (mm_interconnect_0_jtag_avalon_jtag_slave_write),       //                                .write
		.jtag_avalon_jtag_slave_read           (mm_interconnect_0_jtag_avalon_jtag_slave_read),        //                                .read
		.jtag_avalon_jtag_slave_readdata       (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                                .readdata
		.jtag_avalon_jtag_slave_writedata      (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                                .writedata
		.jtag_avalon_jtag_slave_waitrequest    (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.jtag_avalon_jtag_slave_chipselect     (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  //                                .chipselect
		.memory_s1_address                     (mm_interconnect_0_memory_s1_address),                  //                       memory_s1.address
		.memory_s1_write                       (mm_interconnect_0_memory_s1_write),                    //                                .write
		.memory_s1_readdata                    (mm_interconnect_0_memory_s1_readdata),                 //                                .readdata
		.memory_s1_writedata                   (mm_interconnect_0_memory_s1_writedata),                //                                .writedata
		.memory_s1_byteenable                  (mm_interconnect_0_memory_s1_byteenable),               //                                .byteenable
		.memory_s1_chipselect                  (mm_interconnect_0_memory_s1_chipselect),               //                                .chipselect
		.memory_s1_clken                       (mm_interconnect_0_memory_s1_clken),                    //                                .clken
		.out0_s1_address                       (mm_interconnect_0_out0_s1_address),                    //                         out0_s1.address
		.out0_s1_write                         (mm_interconnect_0_out0_s1_write),                      //                                .write
		.out0_s1_readdata                      (mm_interconnect_0_out0_s1_readdata),                   //                                .readdata
		.out0_s1_writedata                     (mm_interconnect_0_out0_s1_writedata),                  //                                .writedata
		.out0_s1_chipselect                    (mm_interconnect_0_out0_s1_chipselect),                 //                                .chipselect
		.out1_s1_address                       (mm_interconnect_0_out1_s1_address),                    //                         out1_s1.address
		.out1_s1_write                         (mm_interconnect_0_out1_s1_write),                      //                                .write
		.out1_s1_readdata                      (mm_interconnect_0_out1_s1_readdata),                   //                                .readdata
		.out1_s1_writedata                     (mm_interconnect_0_out1_s1_writedata),                  //                                .writedata
		.out1_s1_chipselect                    (mm_interconnect_0_out1_s1_chipselect),                 //                                .chipselect
		.out2_s1_address                       (mm_interconnect_0_out2_s1_address),                    //                         out2_s1.address
		.out2_s1_write                         (mm_interconnect_0_out2_s1_write),                      //                                .write
		.out2_s1_readdata                      (mm_interconnect_0_out2_s1_readdata),                   //                                .readdata
		.out2_s1_writedata                     (mm_interconnect_0_out2_s1_writedata),                  //                                .writedata
		.out2_s1_chipselect                    (mm_interconnect_0_out2_s1_chipselect),                 //                                .chipselect
		.out3_s1_address                       (mm_interconnect_0_out3_s1_address),                    //                         out3_s1.address
		.out3_s1_write                         (mm_interconnect_0_out3_s1_write),                      //                                .write
		.out3_s1_readdata                      (mm_interconnect_0_out3_s1_readdata),                   //                                .readdata
		.out3_s1_writedata                     (mm_interconnect_0_out3_s1_writedata),                  //                                .writedata
		.out3_s1_chipselect                    (mm_interconnect_0_out3_s1_chipselect),                 //                                .chipselect
		.out4_s1_address                       (mm_interconnect_0_out4_s1_address),                    //                         out4_s1.address
		.out4_s1_write                         (mm_interconnect_0_out4_s1_write),                      //                                .write
		.out4_s1_readdata                      (mm_interconnect_0_out4_s1_readdata),                   //                                .readdata
		.out4_s1_writedata                     (mm_interconnect_0_out4_s1_writedata),                  //                                .writedata
		.out4_s1_chipselect                    (mm_interconnect_0_out4_s1_chipselect),                 //                                .chipselect
		.out5_s1_address                       (mm_interconnect_0_out5_s1_address),                    //                         out5_s1.address
		.out5_s1_write                         (mm_interconnect_0_out5_s1_write),                      //                                .write
		.out5_s1_readdata                      (mm_interconnect_0_out5_s1_readdata),                   //                                .readdata
		.out5_s1_writedata                     (mm_interconnect_0_out5_s1_writedata),                  //                                .writedata
		.out5_s1_chipselect                    (mm_interconnect_0_out5_s1_chipselect),                 //                                .chipselect
		.out6_s1_address                       (mm_interconnect_0_out6_s1_address),                    //                         out6_s1.address
		.out6_s1_write                         (mm_interconnect_0_out6_s1_write),                      //                                .write
		.out6_s1_readdata                      (mm_interconnect_0_out6_s1_readdata),                   //                                .readdata
		.out6_s1_writedata                     (mm_interconnect_0_out6_s1_writedata),                  //                                .writedata
		.out6_s1_chipselect                    (mm_interconnect_0_out6_s1_chipselect),                 //                                .chipselect
		.out7_s1_address                       (mm_interconnect_0_out7_s1_address),                    //                         out7_s1.address
		.out7_s1_write                         (mm_interconnect_0_out7_s1_write),                      //                                .write
		.out7_s1_readdata                      (mm_interconnect_0_out7_s1_readdata),                   //                                .readdata
		.out7_s1_writedata                     (mm_interconnect_0_out7_s1_writedata),                  //                                .writedata
		.out7_s1_chipselect                    (mm_interconnect_0_out7_s1_chipselect),                 //                                .chipselect
		.out_aux_s1_address                    (mm_interconnect_0_out_aux_s1_address),                 //                      out_aux_s1.address
		.out_aux_s1_write                      (mm_interconnect_0_out_aux_s1_write),                   //                                .write
		.out_aux_s1_readdata                   (mm_interconnect_0_out_aux_s1_readdata),                //                                .readdata
		.out_aux_s1_writedata                  (mm_interconnect_0_out_aux_s1_writedata),               //                                .writedata
		.out_aux_s1_chipselect                 (mm_interconnect_0_out_aux_s1_chipselect),              //                                .chipselect
		.sysid_control_slave_address           (mm_interconnect_0_sysid_control_slave_address),        //             sysid_control_slave.address
		.sysid_control_slave_readdata          (mm_interconnect_0_sysid_control_slave_readdata),       //                                .readdata
		.timer_s1_address                      (mm_interconnect_0_timer_s1_address),                   //                        timer_s1.address
		.timer_s1_write                        (mm_interconnect_0_timer_s1_write),                     //                                .write
		.timer_s1_readdata                     (mm_interconnect_0_timer_s1_readdata),                  //                                .readdata
		.timer_s1_writedata                    (mm_interconnect_0_timer_s1_writedata),                 //                                .writedata
		.timer_s1_chipselect                   (mm_interconnect_0_timer_s1_chipselect)                 //                                .chipselect
	);

	sopc4_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
